module cmd_queue#(parameter DEPTH =16) (

) ; 
// contains fifo



endmodule 