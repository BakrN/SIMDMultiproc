module pool; 


endmodule