`include "proc.sv"
module proc_tb; 


endmodule