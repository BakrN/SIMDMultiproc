// Command Issue
// cores send request here  or could poll 
// contains scoreboard 
module issuer () ; 


endmodule ; 