// Write a test bench 