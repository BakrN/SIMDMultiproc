// Reorder buffer to with CAM containing the cmd_id and proc_ids fields 

module rob ( )